package axiom_apb_pkg;

    `include "config/apb_types.svh"
    `include "config/apb_config.svh"

    `include "seq_items/apb_txn.svh"

    `include "agent/apb_sequencer.svh"
    `include "agent/apb_driver.svh"
    `include "agent/apb_monitor.svh"
    `include "agent/apb_agent.svh"

endpackage
