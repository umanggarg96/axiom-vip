package test_pkg;

    import uvm_pkg::*;
    import axiom_apb_pkg::*;

    `include "uvm_macros.svh"

    `include "env/env.svh"
    `include "env/test_base.svh"

endpackage
