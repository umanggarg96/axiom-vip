typedef enum {
    APB3,
    APB4
} apb_version_t;

typedef enum {
    APB_MASTER,
    APB_SLAVE,
    APB_MONITOR
} apb_agent_t;

